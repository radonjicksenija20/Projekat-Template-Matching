`ifndef CONFIGURATION2_PKG_SV
 `define CONFIGURATION2_PKG_SV

package configurations2_pkg;

   import uvm_pkg::*;      // import the UVM library   
 `include "uvm_macros.svh" // Include the UVM macros

`include "cross_corr_config2.sv"


endpackage : configurations2_pkg

`endif

