`ifndef TEST_BASE_SV
`define TEST_BASE_SV

class test_base extends uvm_test;

   env cross_env;
   cross_corr_config cfg;

   `uvm_component_utils(test_base)

   function new(string name = "test_base", uvm_component parent = null);
      super.new(name,parent);
   endfunction : new

   function void build_phase(uvm_phase phase);
      super.build_phase(phase);
      cfg = cross_corr_config::type_id::create("cfg"); 
      cfg.randomize(); 
      cfg.randomize_config(); //randomize files
      uvm_config_db#(cross_corr_config)::set(this, "cross_env", "cross_corr_config", cfg);      
      cross_env = env::type_id::create("cross_env", this);      
   endfunction : build_phase

   function void end_of_elaboration_phase(uvm_phase phase);
      super.end_of_elaboration_phase(phase);
      uvm_top.print_topology();
   endfunction : end_of_elaboration_phase

endclass : test_base

`endif

